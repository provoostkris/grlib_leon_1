-------------------------------------------------------------------------------
--
-- ROM core VHDL template. See the macro description included
-- behind this frame.
--
-- Copyright (C) 2000 Rudolf Matousek <matousek@utia.cas.cz>
--
-- This code may be used under the terms of Version 2 of the GPL,
-- read the file COPYING for details.
--
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity ROM is
    port(
      clk : in std_logic;
      csn : in std_logic;
      addr : in std_logic_vector (29 downto 0);
      data : out std_logic_vector (31 downto 0)
      );
end ROM;

architecture rtl of ROM is
  signal raddr : std_logic_vector(7 downto 0);
  signal d : std_logic_vector(31 downto 0);
  attribute syn_romstyle : string;
  attribute syn_romstyle of d : signal is "select_rom";
  
begin

  p : process(raddr)
  begin
    case raddr is
    when "00000000" => d <= "10000010000100000010000000000010";
    when "00000001" => d <= "10000001100100000100000000000000";
    when "00000010" => d <= "00000011000000000000000000000100";
    when "00000011" => d <= "10000010000100000110000011000000";
    when "00000100" => d <= "10000001100010000110000000100000";
    when "00000101" => d <= "00000001000000000000000000000000";
    when "00000110" => d <= "00000001000000000000000000000000";
    when "00000111" => d <= "00000001000000000000000000000000";
    when "00001000" => d <= "00000011000000000000000000000000";
    when "00001001" => d <= "10000010000100000110001011111000";
    when "00001010" => d <= "11011100000000000100000000000000";
    when "00001011" => d <= "00000011001000000000000000000000";
    when "00001100" => d <= "11000010000000000110000000010100";
    when "00001101" => d <= "01000000000000000000000010011010";
    when "00001110" => d <= "10011100001000111010000001000000";
    when "00001111" => d <= "10010001110100000010000000000000";
    when "00010000" => d <= "11000110000010100000000000000000";
    when "00010001" => d <= "10000000101000001110000000000000";
    when "00010010" => d <= "00000010100000000000000000001100";
    when "00010011" => d <= "00010011001000000000000000000000";
    when "00010100" => d <= "11000100000000100110000001110100";
    when "00010101" => d <= "10000000100010001010000000000100";
    when "00010110" => d <= "00000010101111111111111111111110";
    when "00010111" => d <= "10000100000010001110000011111111";
    when "00011000" => d <= "11000100001000100110000001110000";
    when "00011001" => d <= "10010000000000100010000000000001";
    when "00011010" => d <= "11000110000010100000000000000000";
    when "00011011" => d <= "10000000101000001110000000000000";
    when "00011100" => d <= "00010010101111111111111111111000";
    when "00011101" => d <= "00000001000000000000000000000000";
    when "00011110" => d <= "10000001110000111110000000001000";
    when "00011111" => d <= "00000001000000000000000000000000";
    when "00100000" => d <= "00010011001000000000000000000000";
    when "00100001" => d <= "11000100000000100110000001110100";
    when "00100010" => d <= "10000000100010001010000000000001";
    when "00100011" => d <= "00000010101111111111111111111110";
    when "00100100" => d <= "00000001000000000000000000000000";
    when "00100101" => d <= "11000100000000100110000001110000";
    when "00100110" => d <= "10000110000010001010000011111111";
    when "00100111" => d <= "10000000101000001110000000001101";
    when "00101000" => d <= "00000010100000000000000000000101";
    when "00101001" => d <= "11000100001010100000000000000000";
    when "00101010" => d <= "10000000101000001110000000001010";
    when "00101011" => d <= "00110010101111111111111111110110";
    when "00101100" => d <= "10010000000000100010000000000001";
    when "00101101" => d <= "10000001110000111110000000001000";
    when "00101110" => d <= "00000001000000000000000000000000";
    when "00101111" => d <= "10010110000100000000000000001000";
    when "00110000" => d <= "10010000000100000010000000000000";
    when "00110001" => d <= "10000000101000100000000000001011";
    when "00110010" => d <= "00010110100000000000000000001101";
    when "00110011" => d <= "10010100000100000010000000000000";
    when "00110100" => d <= "11000100000010100100000000001010";
    when "00110101" => d <= "10000000101000001010000001000000";
    when "00110110" => d <= "00101000100000000000000000000011";
    when "00110111" => d <= "10000100000000001011111111010000";
    when "00111000" => d <= "10000100000000001011111111001001";
    when "00111001" => d <= "10000111001010100010000000000100";
    when "00111010" => d <= "10000100000010001010000011111111";
    when "00111011" => d <= "10010100000000101010000000000001";
    when "00111100" => d <= "10000000101000101000000000001011";
    when "00111101" => d <= "00000110101111111111111111110111";
    when "00111110" => d <= "10010000000100001100000000000010";
    when "00111111" => d <= "10000001110000111110000000001000";
    when "01000000" => d <= "00000001000000000000000000000000";
    when "01000001" => d <= "10011101111000111011111110011000";
    when "01000010" => d <= "10010000000100000010000000000011";
    when "01000011" => d <= "11010000001001100110000000001000";
    when "01000100" => d <= "11010010000011100010000000000001";
    when "01000101" => d <= "10010000000000100111111111001111";
    when "01000110" => d <= "10010000000010100010000011111111";
    when "01000111" => d <= "10000000101000100010000000000010";
    when "01001000" => d <= "00011000100000000000000000001010";
    when "01001001" => d <= "10100000000100000010000000000000";
    when "01001010" => d <= "10010000000100000010000000000001";
    when "01001011" => d <= "01111111111111111111111111100100";
    when "01001100" => d <= "10010010000001100010000000000001";
    when "01001101" => d <= "10010000000000100010000000000001";
    when "01001110" => d <= "10010010000100000010000000000001";
    when "01001111" => d <= "10100001001010100010000000000001";
    when "01010000" => d <= "00010000100000000000000000010101";
    when "01010001" => d <= "11010010001001100110000000001000";
    when "01010010" => d <= "10010000000000100111111111001001";
    when "01010011" => d <= "10010000000010100010000011111111";
    when "01010100" => d <= "10000000101000100010000000000010";
    when "01010101" => d <= "00011000100000000000000000001010";
    when "01010110" => d <= "10010000000100000010000000000001";
    when "01010111" => d <= "01111111111111111111111111011000";
    when "01011000" => d <= "10010010000001100010000000000001";
    when "01011001" => d <= "10010100000100000010000000001011";
    when "01011010" => d <= "10010100001000101000000000001000";
    when "01011011" => d <= "10010010000100000010000000000010";
    when "01011100" => d <= "10100001001010101010000000000001";
    when "01011101" => d <= "00010000100000000000000000001000";
    when "01011110" => d <= "11010010001001100110000000001000";
    when "01011111" => d <= "10010000000010100110000011111111";
    when "01100000" => d <= "10000000101000100010000000110000";
    when "01100001" => d <= "00010010100000000000000000000101";
    when "01100010" => d <= "10010000000100000000000000010000";
    when "01100011" => d <= "10100000000100000010000000000100";
    when "01100100" => d <= "11000000001001100110000000001000";
    when "01100101" => d <= "10010000000100000000000000010000";
    when "01100110" => d <= "01111111111111111111111111001001";
    when "01100111" => d <= "10010010000001100010000000000100";
    when "01101000" => d <= "11010000001001100100000000000000";
    when "01101001" => d <= "10010000000100000010000000000010";
    when "01101010" => d <= "01111111111111111111111111000101";
    when "01101011" => d <= "10010010000001100010000000000010";
    when "01101100" => d <= "10010001001010100010000000000001";
    when "01101101" => d <= "10010000001000100000000000010000";
    when "01101110" => d <= "10010010000001000010000000000100";
    when "01101111" => d <= "10010010000001100000000000001001";
    when "01110000" => d <= "10010000000000100011111111111110";
    when "01110001" => d <= "11010010001001100110000000001100";
    when "01110010" => d <= "11010000001001100110000000000100";
    when "01110011" => d <= "10000001110001111110000000001000";
    when "01110100" => d <= "10000001111010000000000000000000";
    when "01110101" => d <= "00000000000000000000000000000001";
    when "01110110" => d <= "01110011011101000110000101110010";
    when "01110111" => d <= "01110100011010010110111001100111";
    when "01111000" => d <= "00100000011100000111001001101111";
    when "01111001" => d <= "01100111011100100110000101101101";
    when "01111010" => d <= "00111010001000000000101000000000";
    when "01111011" => d <= "10011101111000111011111110011000";
    when "01111100" => d <= "11010000000001100010000000001000";
    when "01111101" => d <= "10000000101000100010000000000001";
    when "01111110" => d <= "00100010100000000000000000000111";
    when "01111111" => d <= "11010000000001100010000000000100";
    when "10000000" => d <= "00001010100000000000000000011101";
    when "10000001" => d <= "10000000101000100010000000000010";
    when "10000010" => d <= "00100010100000000000000000010110";
    when "10000011" => d <= "11100000000001100000000000000000";
    when "10000100" => d <= "00110000100000000000000000011001";
    when "10000101" => d <= "10100000000100000010000000000000";
    when "10000110" => d <= "10010001001100100010000000000001";
    when "10000111" => d <= "10000000101001000000000000001000";
    when "10001000" => d <= "00011010100000000000000000010101";
    when "10001001" => d <= "00000001000000000000000000000000";
    when "10001010" => d <= "11010100000001100010000000001100";
    when "10001011" => d <= "10010011001011000010000000000001";
    when "10001100" => d <= "10010010000000101000000000001001";
    when "10001101" => d <= "01111111111111111111111110100010";
    when "10001110" => d <= "10010000000100000010000000000010";
    when "10001111" => d <= "11010100000001100000000000000000";
    when "10010000" => d <= "11010000001010101000000000010000";
    when "10010001" => d <= "11010010000001100010000000000100";
    when "10010010" => d <= "10100000000001000010000000000001";
    when "10010011" => d <= "10010011001100100110000000000001";
    when "10010100" => d <= "10000000101001000000000000001001";
    when "10010101" => d <= "00101010101111111111111111110110";
    when "10010110" => d <= "11010100000001100010000000001100";
    when "10010111" => d <= "00110000100000000000000000000110";
    when "10011000" => d <= "00010001000000000000000000000000";
    when "10011001" => d <= "01111111111111111111111101110111";
    when "10011010" => d <= "10010000000100100010000111011000";
    when "10011011" => d <= "10011111110001000000000000000000";
    when "10011100" => d <= "00000001000000000000000000000000";
    when "10011101" => d <= "10000001110001111110000000001000";
    when "10011110" => d <= "10000001111010000000000000000000";
    when "10011111" => d <= "00000000000000000000000000000001";
    when "10100000" => d <= "01001100010001010100111101001110";
    when "10100001" => d <= "00100000010100110010110101010010";
    when "10100010" => d <= "01100101011000110110111101110010";
    when "10100011" => d <= "01100100001000000110110001101111";
    when "10100100" => d <= "01100001011001000110010101110010";
    when "10100101" => d <= "00001010000010100000110100111110";
    when "10100110" => d <= "00100000000000000000000000000000";
    when "10100111" => d <= "10011101111000111011111010000000";
    when "10101000" => d <= "01000000000000000000000000010111";
    when "10101001" => d <= "00000001000000000000000000000000";
    when "10101010" => d <= "00010001000000000000000000000000";
    when "10101011" => d <= "01111111111111111111111101100101";
    when "10101100" => d <= "10010000000100100010001010000000";
    when "10101101" => d <= "10100010000001111011111011111000";
    when "10101110" => d <= "10100000000001111011111011100000";
    when "10101111" => d <= "01111111111111111111111101110001";
    when "10110000" => d <= "10010000000100000000000000010001";
    when "10110001" => d <= "11010100000011111011111011111000";
    when "10110010" => d <= "10010000000100000000000000010001";
    when "10110011" => d <= "10000000101000101010000001010011";
    when "10110100" => d <= "00000010100000000000000000000101";
    when "10110101" => d <= "10010010000100000000000000010000";
    when "10110110" => d <= "10000000101000101010000001110011";
    when "10110111" => d <= "00010010101111111111111111111000";
    when "10111000" => d <= "00000001000000000000000000000000";
    when "10111001" => d <= "01111111111111111111111110001000";
    when "10111010" => d <= "00000001000000000000000000000000";
    when "10111011" => d <= "01111111111111111111111111000000";
    when "10111100" => d <= "10010000000100000000000000010000";
    when "10111101" => d <= "00110000101111111111111111110010";
    when "10111110" => d <= "01000000001111111111111111110000";
    when "10111111" => d <= "00010001001000000000000000000000";
    when "11000000" => d <= "11000100000000100010000000010100";
    when "11000001" => d <= "10000000100010001010000000000011";
    when "11000010" => d <= "00010010100000000000000000000111";
    when "11000011" => d <= "00000101000000000000000000101010";
    when "11000100" => d <= "10000001110110000010000000000000";
    when "11000101" => d <= "00000101000000000000000001000000";
    when "11000110" => d <= "10000100000100001010000000001111";
    when "11000111" => d <= "11000100001000100010000000010100";
    when "11001000" => d <= "00000101000000000000000000101010";
    when "11001001" => d <= "10000100000100001010001000000000";
    when "11001010" => d <= "11000100001000100010000010100100";
    when "11001011" => d <= "11000000001000100010000010010000";
    when "11001100" => d <= "11000000001000100010000010010100";
    when "11001101" => d <= "11000000001000100010000010011000";
    when "11001110" => d <= "10000100000100000011111111111111";
    when "11001111" => d <= "11000100001000100010000001000100";
    when "11010000" => d <= "10000110000100000010000000000111";
    when "11010001" => d <= "11000110001000100010000001001000";
    when "11010010" => d <= "11000000001000100010000001110100";
    when "11010011" => d <= "11000000001000100010000010000100";
    when "11010100" => d <= "10000100000100000010000000000011";
    when "11010101" => d <= "11000100001000100010000001111000";
    when "11010110" => d <= "11000100001000100010000010001000";
    when "11010111" => d <= "10000001110000111110000000001000";
    when "11011000" => d <= "00000001000000000000000000000000";
    when "11011001" => d <= "00000000000000000000000000000001";
    when "11011010" => d <= "00000000000000000000000000000001";
    when "11011011" => d <= "00000000000000000000000000000001";

    when others => d <= (others => '-');
    end case;
  end process;

  r : process (clk)
  begin
    if rising_edge(clk) then
      if csn = '0' then raddr <= addr(7 downto 0); end if;
    end if;
  end process;

  data <= d;
end rtl;
